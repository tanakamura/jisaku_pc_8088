parameter AXI_ADDR32_UART_RX = 32'h0x0000000;
parameter AXI_ADDR32_UART_TX = 32'h00000004;
parameter AXI_ADDR32_DRAM_BASE = 32'h80000000;

parameter ADDR_TYPE_INTERNAL_ROM = 3'b000;
parameter ADDR_TYPE_INTERNAL_RAM = 3'b001;
parameter ADDR_TYPE_INTERNAL_LED = 3'b010;
parameter ADDR_TYPE_AXI = 3'b011;
parameter ADDR_TYPE_UNKNOWN = 3'b100;
parameter ADDR_TYPE_NOT_OP = 3'b101;


