parameter AXI_ADDR32_UART_RX = 32'h4060_0000;
parameter AXI_ADDR32_UART_TX = 32'h4060_0004;
parameter AXI_ADDR32_UART_STAT = 32'h4060_0008;
parameter AXI_ADDR32_DRAM_BASE = 32'h8000_0000;
parameter AXI_ADDR32_SPI_FLASH_BASE = 32'h44a0_0000;
parameter AXI_ADDR32_SPI_BASE = 32'h44a1_0000;
parameter AXI_ADDR32_FLASH_XIP_BASE = 32'h0100_0000;

parameter integer ADDR_TYPE_NBIT = 3;

parameter ADDR_TYPE_INTERNAL_ROM = 3'd0;
parameter ADDR_TYPE_INTERNAL_RAM = 3'd1;
parameter ADDR_TYPE_INTERNAL_PERIPHERAL = 3'd2;
parameter ADDR_TYPE_AXI = 3'd5;
parameter ADDR_TYPE_UNKNOWN = 3'd6;
parameter ADDR_TYPE_NOT_OP = 3'd7;


